library ieee;
use ieee.std_logic_1164.all;

entity digital_filter_tb is
end digital_filter_tb;

architecture beh of digital_filter_tb is

component digital_filter is
port ( start : in std_logic;
clock_50,rst : in std_logic;
data_in1: in std_logic_vector(7 downto 0);
done : out std_logic);
end component;
signal start_tb, clk_tb, rst_tb, done_tb: std_logic;
signal input_tb: std_logic_vector(7 downto 0);
begin

testbench: digital_filter port map(start_tb, clk_tb, rst_tb, input_tb, done_tb);
rst_tb <= '0';

clock: process
begin
clk_tb <= '0';
wait for 10 ns;
clk_tb <= '1';
wait for 10 ns;
end process;

segnali: process
begin
input_tb <= "01110001";
start_tb <= '1';
wait for 5 ns;
start_tb <= '0';
wait for 20 ns;
input_tb <= "11001000";
wait for 20 ns;
input_tb <= "10010011";
wait for 20 ns;
input_tb <= "00110011";
wait for 20 ns;
input_tb <= "11111111";
wait for 20 ns;
input_tb <= "10000100";
wait for 20 ns;
input_tb <= "01100111";
wait for 20 ns;
input_tb <= "11011100";
wait for 20 ns;
input_tb <= "11010010";
wait for 20 ns;
input_tb <= "11100110";
wait for 20 ns;
input_tb <= "11110111";
wait for 20 ns;
input_tb <= "01001101";
wait for 20 ns;
input_tb <= "01100000";
wait for 20 ns;
input_tb <= "11010100";
wait for 20 ns;
input_tb <= "10011110";
wait for 20 ns;
input_tb <= "00111111";
wait for 20 ns;
input_tb <= "00010010";
wait for 20 ns;
input_tb <= "01101010";
wait for 20 ns;
input_tb <= "00011011";
wait for 20 ns;
input_tb <= "01001001";
wait for 20 ns;
input_tb <= "10101111";
wait for 20 ns;
input_tb <= "10011101";
wait for 20 ns;
input_tb <= "10011111";
wait for 20 ns;
input_tb <= "10100110";
wait for 20 ns;
input_tb <= "00011000";
wait for 20 ns;
input_tb <= "00011110";
wait for 20 ns;
input_tb <= "00100101";
wait for 20 ns;
input_tb <= "00111001";
wait for 20 ns;
input_tb <= "00110111";
wait for 20 ns;
input_tb <= "10000001";
wait for 20 ns;
input_tb <= "00000010";
wait for 20 ns;
input_tb <= "11001110";
wait for 20 ns;
input_tb <= "00110010";
wait for 20 ns;
input_tb <= "10011111";
wait for 20 ns;
input_tb <= "10111101";
wait for 20 ns;
input_tb <= "10100011";
wait for 20 ns;
input_tb <= "11100100";
wait for 20 ns;
input_tb <= "00111001";
wait for 20 ns;
input_tb <= "00100000";
wait for 20 ns;
input_tb <= "00100111";
wait for 20 ns;
input_tb <= "10001101";
wait for 20 ns;
input_tb <= "11011110";
wait for 20 ns;
input_tb <= "10001111";
wait for 20 ns;
input_tb <= "00000001";
wait for 20 ns;
input_tb <= "11001000";
wait for 20 ns;
input_tb <= "00001110";
wait for 20 ns;
input_tb <= "10011001";
wait for 20 ns;
input_tb <= "01010100";
wait for 20 ns;
input_tb <= "10111110";
wait for 20 ns;
input_tb <= "10011111";
wait for 20 ns;
input_tb <= "11001101";
wait for 20 ns;
input_tb <= "01000001";
wait for 20 ns;
input_tb <= "10011010";
wait for 20 ns;
input_tb <= "01100000";
wait for 20 ns;
input_tb <= "11001111";
wait for 20 ns;
input_tb <= "10101110";
wait for 20 ns;
input_tb <= "00111101";
wait for 20 ns;
input_tb <= "11111101";
wait for 20 ns;
input_tb <= "10101011";
wait for 20 ns;
input_tb <= "01000110";
wait for 20 ns;
input_tb <= "00110010";
wait for 20 ns;
input_tb <= "00100010";
wait for 20 ns;
input_tb <= "01101000";
wait for 20 ns;
input_tb <= "11000001";
wait for 20 ns;
input_tb <= "11100100";
wait for 20 ns;
input_tb <= "11100011";
wait for 20 ns;
input_tb <= "11100001";
wait for 20 ns;
input_tb <= "01100110";
wait for 20 ns;
input_tb <= "00001110";
wait for 20 ns;
input_tb <= "01011100";
wait for 20 ns;
input_tb <= "11010000";
wait for 20 ns;
input_tb <= "11001110";
wait for 20 ns;
input_tb <= "01110100";
wait for 20 ns;
input_tb <= "10010100";
wait for 20 ns;
input_tb <= "00101100";
wait for 20 ns;
input_tb <= "11101010";
wait for 20 ns;
input_tb <= "11010001";
wait for 20 ns;
input_tb <= "10101000";
wait for 20 ns;
input_tb <= "10110101";
wait for 20 ns;
input_tb <= "01001000";
wait for 20 ns;
input_tb <= "00010000";
wait for 20 ns;
input_tb <= "00100101";
wait for 20 ns;
input_tb <= "11001101";
wait for 20 ns;
input_tb <= "10010001";
wait for 20 ns;
input_tb <= "10111110";
wait for 20 ns;
input_tb <= "10110101";
wait for 20 ns;
input_tb <= "10001001";
wait for 20 ns;
input_tb <= "01010111";
wait for 20 ns;
input_tb <= "11000000";
wait for 20 ns;
input_tb <= "11111110";
wait for 20 ns;
input_tb <= "00001000";
wait for 20 ns;
input_tb <= "00001101";
wait for 20 ns;
input_tb <= "01000001";
wait for 20 ns;
input_tb <= "11000111";
wait for 20 ns;
input_tb <= "00000011";
wait for 20 ns;
input_tb <= "01010111";
wait for 20 ns;
input_tb <= "11101111";
wait for 20 ns;
input_tb <= "01011100";
wait for 20 ns;
input_tb <= "10100110";
wait for 20 ns;
input_tb <= "10000101";
wait for 20 ns;
input_tb <= "01100111";
wait for 20 ns;
input_tb <= "00110100";
wait for 20 ns;
input_tb <= "10011110";
wait for 20 ns;
input_tb <= "01011001";
wait for 20 ns;
input_tb <= "11101101";
wait for 20 ns;
input_tb <= "11010010";
wait for 20 ns;
input_tb <= "01110100";
wait for 20 ns;
input_tb <= "00010001";
wait for 20 ns;
input_tb <= "01100001";
wait for 20 ns;
input_tb <= "11101001";
wait for 20 ns;
input_tb <= "00011001";
wait for 20 ns;
input_tb <= "10100001";
wait for 20 ns;
input_tb <= "01101110";
wait for 20 ns;
input_tb <= "11000011";
wait for 20 ns;
input_tb <= "11000010";
wait for 20 ns;
input_tb <= "01000001";
wait for 20 ns;
input_tb <= "00000101";
wait for 20 ns;
input_tb <= "11100011";
wait for 20 ns;
input_tb <= "11110101";
wait for 20 ns;
input_tb <= "00100111";
wait for 20 ns;
input_tb <= "00001010";
wait for 20 ns;
input_tb <= "11101010";
wait for 20 ns;
input_tb <= "11100100";
wait for 20 ns;
input_tb <= "10010110";
wait for 20 ns;
input_tb <= "01001101";
wait for 20 ns;
input_tb <= "10110111";
wait for 20 ns;
input_tb <= "11111011";
wait for 20 ns;
input_tb <= "00010111";
wait for 20 ns;
input_tb <= "10111011";
wait for 20 ns;
input_tb <= "11010010";
wait for 20 ns;
input_tb <= "10110101";
wait for 20 ns;
input_tb <= "00000111";
wait for 20 ns;
input_tb <= "11010110";
wait for 20 ns;
input_tb <= "00001011";
wait for 20 ns;
input_tb <= "10110011";
wait for 20 ns;
input_tb <= "01010001";
wait for 20 ns;
input_tb <= "01100010";
wait for 20 ns;
input_tb <= "01011110";
wait for 20 ns;
input_tb <= "00001111";
wait for 20 ns;
input_tb <= "01111101";
wait for 20 ns;
input_tb <= "01100001";
wait for 20 ns;
input_tb <= "00011010";
wait for 20 ns;
input_tb <= "11101110";
wait for 20 ns;
input_tb <= "11101010";
wait for 20 ns;
input_tb <= "01000010";
wait for 20 ns;
input_tb <= "01000011";
wait for 20 ns;
input_tb <= "01010100";
wait for 20 ns;
input_tb <= "01010111";
wait for 20 ns;
input_tb <= "01010110";
wait for 20 ns;
input_tb <= "00110100";
wait for 20 ns;
input_tb <= "00111101";
wait for 20 ns;
input_tb <= "10101000";
wait for 20 ns;
input_tb <= "10000011";
wait for 20 ns;
input_tb <= "10001000";
wait for 20 ns;
input_tb <= "11101001";
wait for 20 ns;
input_tb <= "11100111";
wait for 20 ns;
input_tb <= "00111100";
wait for 20 ns;
input_tb <= "00111011";
wait for 20 ns;
input_tb <= "01110111";
wait for 20 ns;
input_tb <= "10001010";
wait for 20 ns;
input_tb <= "10110000";
wait for 20 ns;
input_tb <= "00001101";
wait for 20 ns;
input_tb <= "10110101";
wait for 20 ns;
input_tb <= "11110100";
wait for 20 ns;
input_tb <= "01000010";
wait for 20 ns;
input_tb <= "00100111";
wait for 20 ns;
input_tb <= "00110111";
wait for 20 ns;
input_tb <= "00111110";
wait for 20 ns;
input_tb <= "00111010";
wait for 20 ns;
input_tb <= "00000001";
wait for 20 ns;
input_tb <= "10100110";
wait for 20 ns;
input_tb <= "00110110";
wait for 20 ns;
input_tb <= "10111010";
wait for 20 ns;
input_tb <= "10000011";
wait for 20 ns;
input_tb <= "01011011";
wait for 20 ns;
input_tb <= "10101000";
wait for 20 ns;
input_tb <= "11110011";
wait for 20 ns;
input_tb <= "01101011";
wait for 20 ns;
input_tb <= "00101100";
wait for 20 ns;
input_tb <= "11011101";
wait for 20 ns;
input_tb <= "10011000";
wait for 20 ns;
input_tb <= "11101110";
wait for 20 ns;
input_tb <= "10000110";
wait for 20 ns;
input_tb <= "01100010";
wait for 20 ns;
input_tb <= "10010011";
wait for 20 ns;
input_tb <= "10100010";
wait for 20 ns;
input_tb <= "10111101";
wait for 20 ns;
input_tb <= "00001010";
wait for 20 ns;
input_tb <= "11111000";
wait for 20 ns;
input_tb <= "10011011";
wait for 20 ns;
input_tb <= "10011111";
wait for 20 ns;
input_tb <= "00110110";
wait for 20 ns;
input_tb <= "00110111";
wait for 20 ns;
input_tb <= "11010100";
wait for 20 ns;
input_tb <= "01001111";
wait for 20 ns;
input_tb <= "01010100";
wait for 20 ns;
input_tb <= "10010101";
wait for 20 ns;
input_tb <= "11010001";
wait for 20 ns;
input_tb <= "01010001";
wait for 20 ns;
input_tb <= "10100110";
wait for 20 ns;
input_tb <= "11011101";
wait for 20 ns;
input_tb <= "10000011";
wait for 20 ns;
input_tb <= "11100001";
wait for 20 ns;
input_tb <= "01000101";
wait for 20 ns;
input_tb <= "01010010";
wait for 20 ns;
input_tb <= "01101100";
wait for 20 ns;
input_tb <= "10001001";
wait for 20 ns;
input_tb <= "01100101";
wait for 20 ns;
input_tb <= "11101001";
wait for 20 ns;
input_tb <= "00000100";
wait for 20 ns;
input_tb <= "11110010";
wait for 20 ns;
input_tb <= "11011010";
wait for 20 ns;
input_tb <= "10110101";
wait for 20 ns;
input_tb <= "01011010";
wait for 20 ns;
input_tb <= "11111011";
wait for 20 ns;
input_tb <= "11011100";
wait for 20 ns;
input_tb <= "10100011";
wait for 20 ns;
input_tb <= "11111110";
wait for 20 ns;
input_tb <= "00001000";
wait for 20 ns;
input_tb <= "00000111";
wait for 20 ns;
input_tb <= "01100111";
wait for 20 ns;
input_tb <= "00011111";
wait for 20 ns;
input_tb <= "10011100";
wait for 20 ns;
input_tb <= "10100101";
wait for 20 ns;
input_tb <= "10110110";
wait for 20 ns;
input_tb <= "11110001";
wait for 20 ns;
input_tb <= "00101011";
wait for 20 ns;
input_tb <= "00110000";
wait for 20 ns;
input_tb <= "10110110";
wait for 20 ns;
input_tb <= "01010001";
wait for 20 ns;
input_tb <= "00101001";
wait for 20 ns;
input_tb <= "00010011";
wait for 20 ns;
input_tb <= "10110011";
wait for 20 ns;
input_tb <= "10101100";
wait for 20 ns;
input_tb <= "01100111";
wait for 20 ns;
input_tb <= "10110001";
wait for 20 ns;
input_tb <= "00010011";
wait for 20 ns;
input_tb <= "00011101";
wait for 20 ns;
input_tb <= "10011111";
wait for 20 ns;
input_tb <= "10101000";
wait for 20 ns;
input_tb <= "10001100";
wait for 20 ns;
input_tb <= "11010101";
wait for 20 ns;
input_tb <= "01001110";
wait for 20 ns;
input_tb <= "01010111";
wait for 20 ns;
input_tb <= "10010100";
wait for 20 ns;
input_tb <= "11000000";
wait for 20 ns;
input_tb <= "11000001";
wait for 20 ns;
input_tb <= "10011110";
wait for 20 ns;
input_tb <= "00011001";
wait for 20 ns;
input_tb <= "01100110";
wait for 20 ns;
input_tb <= "01110011";
wait for 20 ns;
input_tb <= "11100100";
wait for 20 ns;
input_tb <= "01110011";
wait for 20 ns;
input_tb <= "00001111";
wait for 20 ns;
input_tb <= "10010110";
wait for 20 ns;
input_tb <= "01011111";
wait for 20 ns;
input_tb <= "10010111";
wait for 20 ns;
input_tb <= "00101010";
wait for 20 ns;
input_tb <= "11110000";
wait for 20 ns;
input_tb <= "10001111";
wait for 20 ns;
input_tb <= "10001101";
wait for 20 ns;
input_tb <= "11101111";
wait for 20 ns;
input_tb <= "11101000";
wait for 20 ns;
input_tb <= "00001100";
wait for 20 ns;
input_tb <= "00100100";
wait for 20 ns;
input_tb <= "01000100";
wait for 20 ns;
input_tb <= "11100001";
wait for 20 ns;
input_tb <= "10000010";
wait for 20 ns;
input_tb <= "11100100";
wait for 20 ns;
input_tb <= "11011101";
wait for 20 ns;
input_tb <= "11000110";
wait for 20 ns;
input_tb <= "11111010";
wait for 20 ns;
input_tb <= "01000100";
wait for 20 ns;
input_tb <= "10101000";
wait for 20 ns;
input_tb <= "11100110";
wait for 20 ns;
input_tb <= "01011011";
wait for 20 ns;
input_tb <= "00011101";
wait for 20 ns;
input_tb <= "01101000";
wait for 20 ns;
input_tb <= "00000011";
wait for 20 ns;
input_tb <= "00110000";
wait for 20 ns;
input_tb <= "01011111";
wait for 20 ns;
input_tb <= "10011111";
wait for 20 ns;
input_tb <= "10100101";
wait for 20 ns;
input_tb <= "10101011";
wait for 20 ns;
input_tb <= "00000011";
wait for 20 ns;
input_tb <= "10110010";
wait for 20 ns;
input_tb <= "10110100";
wait for 20 ns;
input_tb <= "11101010";
wait for 20 ns;
input_tb <= "01000000";
wait for 20 ns;
input_tb <= "01001000";
wait for 20 ns;
input_tb <= "01000110";
wait for 20 ns;
input_tb <= "01111010";
wait for 20 ns;
input_tb <= "00000010";
wait for 20 ns;
input_tb <= "11110011";
wait for 20 ns;
input_tb <= "10110110";
wait for 20 ns;
input_tb <= "00011010";
wait for 20 ns;
input_tb <= "10011000";
wait for 20 ns;
input_tb <= "00010010";
wait for 20 ns;
input_tb <= "11110110";
wait for 20 ns;
input_tb <= "11000001";
wait for 20 ns;
input_tb <= "10101100";
wait for 20 ns;
input_tb <= "11110110";
wait for 20 ns;
input_tb <= "00100110";
wait for 20 ns;
input_tb <= "11100010";
wait for 20 ns;
input_tb <= "01111001";
wait for 20 ns;
input_tb <= "01000011";
wait for 20 ns;
input_tb <= "01100101";
wait for 20 ns;
input_tb <= "11101110";
wait for 20 ns;
input_tb <= "00111000";
wait for 20 ns;
input_tb <= "10011001";
wait for 20 ns;
input_tb <= "11100111";
wait for 20 ns;
input_tb <= "00011011";
wait for 20 ns;
input_tb <= "11011011";
wait for 20 ns;
input_tb <= "01110100";
wait for 20 ns;
input_tb <= "01000111";
wait for 20 ns;
input_tb <= "01100100";
wait for 20 ns;
input_tb <= "11111110";
wait for 20 ns;
input_tb <= "01010001";
wait for 20 ns;
input_tb <= "00011111";
wait for 20 ns;
input_tb <= "11010000";
wait for 20 ns;
input_tb <= "00011011";
wait for 20 ns;
input_tb <= "00010011";
wait for 20 ns;
input_tb <= "11010111";
wait for 20 ns;
input_tb <= "11111000";
wait for 20 ns;
input_tb <= "11111101";
wait for 20 ns;
input_tb <= "10100100";
wait for 20 ns;
input_tb <= "10111010";
wait for 20 ns;
input_tb <= "11000011";
wait for 20 ns;
input_tb <= "01110111";
wait for 20 ns;
input_tb <= "11011111";
wait for 20 ns;
input_tb <= "01001111";
wait for 20 ns;
input_tb <= "01110101";
wait for 20 ns;
input_tb <= "01010101";
wait for 20 ns;
input_tb <= "10101110";
wait for 20 ns;
input_tb <= "11100110";
wait for 20 ns;
input_tb <= "11101000";
wait for 20 ns;
input_tb <= "10010011";
wait for 20 ns;
input_tb <= "01101111";
wait for 20 ns;
input_tb <= "01110001";
wait for 20 ns;
input_tb <= "00011000";
wait for 20 ns;
input_tb <= "11001101";
wait for 20 ns;
input_tb <= "10011101";
wait for 20 ns;
input_tb <= "10010101";
wait for 20 ns;
input_tb <= "11100110";
wait for 20 ns;
input_tb <= "11110111";
wait for 20 ns;
input_tb <= "10101100";
wait for 20 ns;
input_tb <= "00000001";
wait for 20 ns;
input_tb <= "00010101";
wait for 20 ns;
input_tb <= "01001110";
wait for 20 ns;
input_tb <= "00110100";
wait for 20 ns;
input_tb <= "11111111";
wait for 20 ns;
input_tb <= "10011001";
wait for 20 ns;
input_tb <= "10001110";
wait for 20 ns;
input_tb <= "01010010";
wait for 20 ns;
input_tb <= "01001000";
wait for 20 ns;
input_tb <= "00010001";
wait for 20 ns;
input_tb <= "01100110";
wait for 20 ns;
input_tb <= "01001100";
wait for 20 ns;
input_tb <= "00011101";
wait for 20 ns;
input_tb <= "10010010";
wait for 20 ns;
input_tb <= "00101001";
wait for 20 ns;
input_tb <= "01110011";
wait for 20 ns;
input_tb <= "10010011";
wait for 20 ns;
input_tb <= "10100110";
wait for 20 ns;
input_tb <= "11000110";
wait for 20 ns;
input_tb <= "01001110";
wait for 20 ns;
input_tb <= "00101111";
wait for 20 ns;
input_tb <= "10010100";
wait for 20 ns;
input_tb <= "11111010";
wait for 20 ns;
input_tb <= "11110100";
wait for 20 ns;
input_tb <= "10110010";
wait for 20 ns;
input_tb <= "11100010";
wait for 20 ns;
input_tb <= "11000100";
wait for 20 ns;
input_tb <= "10111010";
wait for 20 ns;
input_tb <= "00110110";
wait for 20 ns;
input_tb <= "00011001";
wait for 20 ns;
input_tb <= "00011010";
wait for 20 ns;
input_tb <= "00001110";
wait for 20 ns;
input_tb <= "01111010";
wait for 20 ns;
input_tb <= "11001000";
wait for 20 ns;
input_tb <= "11011010";
wait for 20 ns;
input_tb <= "10100011";
wait for 20 ns;
input_tb <= "01111011";
wait for 20 ns;
input_tb <= "11001011";
wait for 20 ns;
input_tb <= "00000011";
wait for 20 ns;
input_tb <= "11001111";
wait for 20 ns;
input_tb <= "01000100";
wait for 20 ns;
input_tb <= "11001101";
wait for 20 ns;
input_tb <= "00100101";
wait for 20 ns;
input_tb <= "00110001";
wait for 20 ns;
input_tb <= "00000110";
wait for 20 ns;
input_tb <= "00001100";
wait for 20 ns;
input_tb <= "00010110";
wait for 20 ns;
input_tb <= "10010110";
wait for 20 ns;
input_tb <= "01101011";
wait for 20 ns;
input_tb <= "01011100";
wait for 20 ns;
input_tb <= "11100111";
wait for 20 ns;
input_tb <= "00011101";
wait for 20 ns;
input_tb <= "00101000";
wait for 20 ns;
input_tb <= "01101111";
wait for 20 ns;
input_tb <= "00010110";
wait for 20 ns;
input_tb <= "10011010";
wait for 20 ns;
input_tb <= "11010010";
wait for 20 ns;
input_tb <= "01010011";
wait for 20 ns;
input_tb <= "00000101";
wait for 20 ns;
input_tb <= "00111001";
wait for 20 ns;
input_tb <= "11110010";
wait for 20 ns;
input_tb <= "00111100";
wait for 20 ns;
input_tb <= "10101011";
wait for 20 ns;
input_tb <= "01100100";
wait for 20 ns;
input_tb <= "01011011";
wait for 20 ns;
input_tb <= "10000100";
wait for 20 ns;
input_tb <= "10001010";
wait for 20 ns;
input_tb <= "11100110";
wait for 20 ns;
input_tb <= "10111011";
wait for 20 ns;
input_tb <= "11110000";
wait for 20 ns;
input_tb <= "11100001";
wait for 20 ns;
input_tb <= "01010000";
wait for 20 ns;
input_tb <= "01110001";
wait for 20 ns;
input_tb <= "00110101";
wait for 20 ns;
input_tb <= "00100010";
wait for 20 ns;
input_tb <= "10011011";
wait for 20 ns;
input_tb <= "10011110";
wait for 20 ns;
input_tb <= "10111011";
wait for 20 ns;
input_tb <= "10100110";
wait for 20 ns;
input_tb <= "00010000";
wait for 20 ns;
input_tb <= "01111111";
wait for 20 ns;
input_tb <= "10100000";
wait for 20 ns;
input_tb <= "10100000";
wait for 20 ns;
input_tb <= "01100101";
wait for 20 ns;
input_tb <= "11111010";
wait for 20 ns;
input_tb <= "00000000";
wait for 20 ns;
input_tb <= "01010000";
wait for 20 ns;
input_tb <= "00101001";
wait for 20 ns;
input_tb <= "01110110";
wait for 20 ns;
input_tb <= "01110100";
wait for 20 ns;
input_tb <= "01111001";
wait for 20 ns;
input_tb <= "01100010";
wait for 20 ns;
input_tb <= "11110000";
wait for 20 ns;
input_tb <= "11011000";
wait for 20 ns;
input_tb <= "00010100";
wait for 20 ns;
input_tb <= "01110100";
wait for 20 ns;
input_tb <= "01001011";
wait for 20 ns;
input_tb <= "01010010";
wait for 20 ns;
input_tb <= "01000110";
wait for 20 ns;
input_tb <= "01000100";
wait for 20 ns;
input_tb <= "11101000";
wait for 20 ns;
input_tb <= "10001111";
wait for 20 ns;
input_tb <= "10010000";
wait for 20 ns;
input_tb <= "10011110";
wait for 20 ns;
input_tb <= "01110111";
wait for 20 ns;
input_tb <= "01010000";
wait for 20 ns;
input_tb <= "01000110";
wait for 20 ns;
input_tb <= "11010100";
wait for 20 ns;
input_tb <= "00001101";
wait for 20 ns;
input_tb <= "00100110";
wait for 20 ns;
input_tb <= "01000010";
wait for 20 ns;
input_tb <= "10101000";
wait for 20 ns;
input_tb <= "01110110";
wait for 20 ns;
input_tb <= "01111001";
wait for 20 ns;
input_tb <= "11011001";
wait for 20 ns;
input_tb <= "01101100";
wait for 20 ns;
input_tb <= "11001100";
wait for 20 ns;
input_tb <= "11001111";
wait for 20 ns;
input_tb <= "00001110";
wait for 20 ns;
input_tb <= "01101000";
wait for 20 ns;
input_tb <= "01001000";
wait for 20 ns;
input_tb <= "01001011";
wait for 20 ns;
input_tb <= "00000110";
wait for 20 ns;
input_tb <= "01111100";
wait for 20 ns;
input_tb <= "01011001";
wait for 20 ns;
input_tb <= "01110100";
wait for 20 ns;
input_tb <= "10111100";
wait for 20 ns;
input_tb <= "00000111";
wait for 20 ns;
input_tb <= "11110011";
wait for 20 ns;
input_tb <= "00111001";
wait for 20 ns;
input_tb <= "11110110";
wait for 20 ns;
input_tb <= "00000111";
wait for 20 ns;
input_tb <= "00101010";
wait for 20 ns;
input_tb <= "00110001";
wait for 20 ns;
input_tb <= "01111000";
wait for 20 ns;
input_tb <= "10000001";
wait for 20 ns;
input_tb <= "11111111";
wait for 20 ns;
input_tb <= "00100111";
wait for 20 ns;
input_tb <= "01110111";
wait for 20 ns;
input_tb <= "00100011";
wait for 20 ns;
input_tb <= "01111010";
wait for 20 ns;
input_tb <= "11010101";
wait for 20 ns;
input_tb <= "01010000";
wait for 20 ns;
input_tb <= "00101000";
wait for 20 ns;
input_tb <= "11111001";
wait for 20 ns;
input_tb <= "11110000";
wait for 20 ns;
input_tb <= "01111010";
wait for 20 ns;
input_tb <= "01111100";
wait for 20 ns;
input_tb <= "11000111";
wait for 20 ns;
input_tb <= "01100101";
wait for 20 ns;
input_tb <= "10111001";
wait for 20 ns;
input_tb <= "00100000";
wait for 20 ns;
input_tb <= "11110000";
wait for 20 ns;
input_tb <= "11100011";
wait for 20 ns;
input_tb <= "10010101";
wait for 20 ns;
input_tb <= "11010001";
wait for 20 ns;
input_tb <= "01010100";
wait for 20 ns;
input_tb <= "10011001";
wait for 20 ns;
input_tb <= "00001011";
wait for 20 ns;
input_tb <= "11100100";
wait for 20 ns;
input_tb <= "11111011";
wait for 20 ns;
input_tb <= "01000001";
wait for 20 ns;
input_tb <= "10000010";
wait for 20 ns;
input_tb <= "01110101";
wait for 20 ns;
input_tb <= "10101000";
wait for 20 ns;
input_tb <= "01011101";
wait for 20 ns;
input_tb <= "00000001";
wait for 20 ns;
input_tb <= "11000000";
wait for 20 ns;
input_tb <= "10110001";
wait for 20 ns;
input_tb <= "11000000";
wait for 20 ns;
input_tb <= "10011110";
wait for 20 ns;
input_tb <= "11001111";
wait for 20 ns;
input_tb <= "00001101";
wait for 20 ns;
input_tb <= "01010001";
wait for 20 ns;
input_tb <= "00111010";
wait for 20 ns;
input_tb <= "01010110";
wait for 20 ns;
input_tb <= "10101111";
wait for 20 ns;
input_tb <= "00001100";
wait for 20 ns;
input_tb <= "01101011";
wait for 20 ns;
input_tb <= "11011011";
wait for 20 ns;
input_tb <= "00010010";
wait for 20 ns;
input_tb <= "01001001";
wait for 20 ns;
input_tb <= "10111010";
wait for 20 ns;
input_tb <= "00011001";
wait for 20 ns;
input_tb <= "00010110";
wait for 20 ns;
input_tb <= "01000001";
wait for 20 ns;
input_tb <= "00001111";
wait for 20 ns;
input_tb <= "10100111";
wait for 20 ns;
input_tb <= "00001010";
wait for 20 ns;
input_tb <= "11001110";
wait for 20 ns;
input_tb <= "01101001";
wait for 20 ns;
input_tb <= "11010101";
wait for 20 ns;
input_tb <= "00001010";
wait for 20 ns;
input_tb <= "01110010";
wait for 20 ns;
input_tb <= "11010010";
wait for 20 ns;
input_tb <= "11010111";
wait for 20 ns;
input_tb <= "10001011";
wait for 20 ns;
input_tb <= "10011011";
wait for 20 ns;
input_tb <= "10010011";
wait for 20 ns;
input_tb <= "00100101";
wait for 20 ns;
input_tb <= "00110100";
wait for 20 ns;
input_tb <= "00100101";
wait for 20 ns;
input_tb <= "10100100";
wait for 20 ns;
input_tb <= "00100001";
wait for 20 ns;
input_tb <= "11110000";
wait for 20 ns;
input_tb <= "00100001";
wait for 20 ns;
input_tb <= "01100110";
wait for 20 ns;
input_tb <= "11111010";
wait for 20 ns;
input_tb <= "01000001";
wait for 20 ns;
input_tb <= "11010101";
wait for 20 ns;
input_tb <= "10010100";
wait for 20 ns;
input_tb <= "11010001";
wait for 20 ns;
input_tb <= "11010111";
wait for 20 ns;
input_tb <= "00000011";
wait for 20 ns;
input_tb <= "01110111";
wait for 20 ns;
input_tb <= "00011011";
wait for 20 ns;
input_tb <= "01100001";
wait for 20 ns;
input_tb <= "01101111";
wait for 20 ns;
input_tb <= "01011010";
wait for 20 ns;
input_tb <= "01000111";
wait for 20 ns;
input_tb <= "10100011";
wait for 20 ns;
input_tb <= "10011011";
wait for 20 ns;
input_tb <= "00111110";
wait for 20 ns;
input_tb <= "10100000";
wait for 20 ns;
input_tb <= "11001000";
wait for 20 ns;
input_tb <= "11010101";
wait for 20 ns;
input_tb <= "11001111";
wait for 20 ns;
input_tb <= "01110100";
wait for 20 ns;
input_tb <= "11111010";
wait for 20 ns;
input_tb <= "01110011";
wait for 20 ns;
input_tb <= "10010110";
wait for 20 ns;
input_tb <= "01110110";
wait for 20 ns;
input_tb <= "00110001";
wait for 20 ns;
input_tb <= "01011110";
wait for 20 ns;
input_tb <= "01101111";
wait for 20 ns;
input_tb <= "01100001";
wait for 20 ns;
input_tb <= "01001000";
wait for 20 ns;
input_tb <= "11001101";
wait for 20 ns;
input_tb <= "00111110";
wait for 20 ns;
input_tb <= "11011110";
wait for 20 ns;
input_tb <= "01010110";
wait for 20 ns;
input_tb <= "01010011";
wait for 20 ns;
input_tb <= "11011110";
wait for 20 ns;
input_tb <= "10101000";
wait for 20 ns;
input_tb <= "00111011";
wait for 20 ns;
input_tb <= "00011100";
wait for 20 ns;
input_tb <= "01011010";
wait for 20 ns;
input_tb <= "11101110";
wait for 20 ns;
input_tb <= "01111001";
wait for 20 ns;
input_tb <= "01110100";
wait for 20 ns;
input_tb <= "01100000";
wait for 20 ns;
input_tb <= "11111001";
wait for 20 ns;
input_tb <= "01000110";
wait for 20 ns;
input_tb <= "10001000";
wait for 20 ns;
input_tb <= "11110010";
wait for 20 ns;
input_tb <= "00001110";
wait for 20 ns;
input_tb <= "11011111";
wait for 20 ns;
input_tb <= "01110001";
wait for 20 ns;
input_tb <= "01011111";
wait for 20 ns;
input_tb <= "10010110";
wait for 20 ns;
input_tb <= "00011110";
wait for 20 ns;
input_tb <= "01101110";
wait for 20 ns;
input_tb <= "01110010";
wait for 20 ns;
input_tb <= "01111100";
wait for 20 ns;
input_tb <= "01001111";
wait for 20 ns;
input_tb <= "01110001";
wait for 20 ns;
input_tb <= "11101001";
wait for 20 ns;
input_tb <= "11010111";
wait for 20 ns;
input_tb <= "01000000";
wait for 20 ns;
input_tb <= "11011110";
wait for 20 ns;
input_tb <= "00101000";
wait for 20 ns;
input_tb <= "11001001";
wait for 20 ns;
input_tb <= "10010111";
wait for 20 ns;
input_tb <= "10001111";
wait for 20 ns;
input_tb <= "00101111";
wait for 20 ns;
input_tb <= "10100110";
wait for 20 ns;
input_tb <= "01101000";
wait for 20 ns;
input_tb <= "00011011";
wait for 20 ns;
input_tb <= "11001010";
wait for 20 ns;
input_tb <= "01011001";
wait for 20 ns;
input_tb <= "00000111";
wait for 20 ns;
input_tb <= "01011000";
wait for 20 ns;
input_tb <= "00000111";
wait for 20 ns;
input_tb <= "00000100";
wait for 20 ns;
input_tb <= "00011011";
wait for 20 ns;
input_tb <= "00011110";
wait for 20 ns;
input_tb <= "11101101";
wait for 20 ns;
input_tb <= "11100111";
wait for 20 ns;
input_tb <= "11110100";
wait for 20 ns;
input_tb <= "01001110";
wait for 20 ns;
input_tb <= "01101011";
wait for 20 ns;
input_tb <= "10000011";
wait for 20 ns;
input_tb <= "00011111";
wait for 20 ns;
input_tb <= "00010011";
wait for 20 ns;
input_tb <= "10001111";
wait for 20 ns;
input_tb <= "11111111";
wait for 20 ns;
input_tb <= "00110111";
wait for 20 ns;
input_tb <= "01101000";
wait for 20 ns;
input_tb <= "11111001";
wait for 20 ns;
input_tb <= "11001010";
wait for 20 ns;
input_tb <= "11111101";
wait for 20 ns;
input_tb <= "11011011";
wait for 20 ns;
input_tb <= "10001110";
wait for 20 ns;
input_tb <= "10000010";
wait for 20 ns;
input_tb <= "10101011";
wait for 20 ns;
input_tb <= "10010000";
wait for 20 ns;
input_tb <= "01110001";
wait for 20 ns;
input_tb <= "00010101";
wait for 20 ns;
input_tb <= "10000110";
wait for 20 ns;
input_tb <= "10001000";
wait for 20 ns;
input_tb <= "00101111";
wait for 20 ns;
input_tb <= "00100110";
wait for 20 ns;
input_tb <= "10110011";
wait for 20 ns;
input_tb <= "00100011";
wait for 20 ns;
input_tb <= "00111001";
wait for 20 ns;
input_tb <= "10110010";
wait for 20 ns;
input_tb <= "01001011";
wait for 20 ns;
input_tb <= "11100100";
wait for 20 ns;
input_tb <= "10011000";
wait for 20 ns;
input_tb <= "11110011";
wait for 20 ns;
input_tb <= "10110010";
wait for 20 ns;
input_tb <= "01110101";
wait for 20 ns;
input_tb <= "11011100";
wait for 20 ns;
input_tb <= "10000100";
wait for 20 ns;
input_tb <= "00100100";
wait for 20 ns;
input_tb <= "11101011";
wait for 20 ns;
input_tb <= "01010101";
wait for 20 ns;
input_tb <= "11000111";
wait for 20 ns;
input_tb <= "10010000";
wait for 20 ns;
input_tb <= "01001010";
wait for 20 ns;
input_tb <= "10000110";
wait for 20 ns;
input_tb <= "10000100";
wait for 20 ns;
input_tb <= "10101010";
wait for 20 ns;
input_tb <= "01001100";
wait for 20 ns;
input_tb <= "11010111";
wait for 20 ns;
input_tb <= "11010010";
wait for 20 ns;
input_tb <= "00111100";
wait for 20 ns;
input_tb <= "01011110";
wait for 20 ns;
input_tb <= "10001010";
wait for 20 ns;
input_tb <= "00111011";
wait for 20 ns;
input_tb <= "10111100";
wait for 20 ns;
input_tb <= "11101100";
wait for 20 ns;
input_tb <= "11110000";
wait for 20 ns;
input_tb <= "00011011";
wait for 20 ns;
input_tb <= "00100100";
wait for 20 ns;
input_tb <= "11011110";
wait for 20 ns;
input_tb <= "11011101";
wait for 20 ns;
input_tb <= "01001001";
wait for 20 ns;
input_tb <= "11111110";
wait for 20 ns;
input_tb <= "01100011";
wait for 20 ns;
input_tb <= "01011001";
wait for 20 ns;
input_tb <= "11111001";
wait for 20 ns;
input_tb <= "10111110";
wait for 20 ns;
input_tb <= "11101101";
wait for 20 ns;
input_tb <= "10011000";
wait for 20 ns;
input_tb <= "11100001";
wait for 20 ns;
input_tb <= "01010101";
wait for 20 ns;
input_tb <= "01111101";
wait for 20 ns;
input_tb <= "00101101";
wait for 20 ns;
input_tb <= "10011011";
wait for 20 ns;
input_tb <= "00000011";
wait for 20 ns;
input_tb <= "00100000";
wait for 20 ns;
input_tb <= "01111010";
wait for 20 ns;
input_tb <= "01001011";
wait for 20 ns;
input_tb <= "01101101";
wait for 20 ns;
input_tb <= "10111001";
wait for 20 ns;
input_tb <= "01101011";
wait for 20 ns;
input_tb <= "10000001";
wait for 20 ns;
input_tb <= "11101111";
wait for 20 ns;
input_tb <= "00000010";
wait for 20 ns;
input_tb <= "01100100";
wait for 20 ns;
input_tb <= "01100001";
wait for 20 ns;
input_tb <= "00110011";
wait for 20 ns;
input_tb <= "11001110";
wait for 20 ns;
input_tb <= "01110111";
wait for 20 ns;
input_tb <= "00000001";
wait for 20 ns;
input_tb <= "00000011";
wait for 20 ns;
input_tb <= "10010001";
wait for 20 ns;
input_tb <= "11011011";
wait for 20 ns;
input_tb <= "00010010";
wait for 20 ns;
input_tb <= "01011011";
wait for 20 ns;
input_tb <= "00100001";
wait for 20 ns;
input_tb <= "10011001";
wait for 20 ns;
input_tb <= "11000011";
wait for 20 ns;
input_tb <= "11000011";
wait for 20 ns;
input_tb <= "10111110";
wait for 20 ns;
input_tb <= "10001001";
wait for 20 ns;
input_tb <= "11100010";
wait for 20 ns;
input_tb <= "11011011";
wait for 20 ns;
input_tb <= "01010001";
wait for 20 ns;
input_tb <= "01111101";
wait for 20 ns;
input_tb <= "01000100";
wait for 20 ns;
input_tb <= "00111000";
wait for 20 ns;
input_tb <= "11110001";
wait for 20 ns;
input_tb <= "10111100";
wait for 20 ns;
input_tb <= "01101000";
wait for 20 ns;
input_tb <= "01101110";
wait for 20 ns;
input_tb <= "10101011";
wait for 20 ns;
input_tb <= "10110010";
wait for 20 ns;
input_tb <= "01010111";
wait for 20 ns;
input_tb <= "01101110";
wait for 20 ns;
input_tb <= "10000011";
wait for 20 ns;
input_tb <= "11100101";
wait for 20 ns;
input_tb <= "11001110";
wait for 20 ns;
input_tb <= "00010011";
wait for 20 ns;
input_tb <= "10110110";
wait for 20 ns;
input_tb <= "00101011";
wait for 20 ns;
input_tb <= "10011111";
wait for 20 ns;
input_tb <= "11110111";
wait for 20 ns;
input_tb <= "01000010";
wait for 20 ns;
input_tb <= "00011011";
wait for 20 ns;
input_tb <= "01010101";
wait for 20 ns;
input_tb <= "10001011";
wait for 20 ns;
input_tb <= "10101000";
wait for 20 ns;
input_tb <= "11000001";
wait for 20 ns;
input_tb <= "00010111";
wait for 20 ns;
input_tb <= "01100111";
wait for 20 ns;
input_tb <= "11110001";
wait for 20 ns;
input_tb <= "10010110";
wait for 20 ns;
input_tb <= "11001111";
wait for 20 ns;
input_tb <= "11011110";
wait for 20 ns;
input_tb <= "11101111";
wait for 20 ns;
input_tb <= "10101110";
wait for 20 ns;
input_tb <= "10001011";
wait for 20 ns;
input_tb <= "11010110";
wait for 20 ns;
input_tb <= "11000101";
wait for 20 ns;
input_tb <= "00110100";
wait for 20 ns;
input_tb <= "00100011";
wait for 20 ns;
input_tb <= "11010110";
wait for 20 ns;
input_tb <= "10101010";
wait for 20 ns;
input_tb <= "00010100";
wait for 20 ns;
input_tb <= "00011100";
wait for 20 ns;
input_tb <= "01100001";
wait for 20 ns;
input_tb <= "11101001";
wait for 20 ns;
input_tb <= "11110111";
wait for 20 ns;
input_tb <= "11001100";
wait for 20 ns;
input_tb <= "10000011";
wait for 20 ns;
input_tb <= "00101100";
wait for 20 ns;
input_tb <= "01110100";
wait for 20 ns;
input_tb <= "10111111";
wait for 20 ns;
input_tb <= "10101001";
wait for 20 ns;
input_tb <= "11111011";
wait for 20 ns;
input_tb <= "10000100";
wait for 20 ns;
input_tb <= "01011010";
wait for 20 ns;
input_tb <= "10110110";
wait for 20 ns;
input_tb <= "10000000";
wait for 20 ns;
input_tb <= "00110111";
wait for 20 ns;
input_tb <= "10111110";
wait for 20 ns;
input_tb <= "01010010";
wait for 20 ns;
input_tb <= "10001101";
wait for 20 ns;
input_tb <= "10100110";
wait for 20 ns;
input_tb <= "11101111";
wait for 20 ns;
input_tb <= "10000101";
wait for 20 ns;
input_tb <= "11100000";
wait for 20 ns;
input_tb <= "00101001";
wait for 20 ns;
input_tb <= "00110110";
wait for 20 ns;
input_tb <= "10000110";
wait for 20 ns;
input_tb <= "10100101";
wait for 20 ns;
input_tb <= "11001010";
wait for 20 ns;
input_tb <= "11000011";
wait for 20 ns;
input_tb <= "11001101";
wait for 20 ns;
input_tb <= "00111100";
wait for 20 ns;
input_tb <= "11111001";
wait for 20 ns;
input_tb <= "10010111";
wait for 20 ns;
input_tb <= "01101111";
wait for 20 ns;
input_tb <= "00111101";
wait for 20 ns;
input_tb <= "10000001";
wait for 20 ns;
input_tb <= "10100001";
wait for 20 ns;
input_tb <= "10101011";
wait for 20 ns;
input_tb <= "10111001";
wait for 20 ns;
input_tb <= "10111010";
wait for 20 ns;
input_tb <= "00100111";
wait for 20 ns;
input_tb <= "11000000";
wait for 20 ns;
input_tb <= "11000011";
wait for 20 ns;
input_tb <= "00000000";
wait for 20 ns;
input_tb <= "01101000";
wait for 20 ns;
input_tb <= "00000010";
wait for 20 ns;
input_tb <= "00101111";
wait for 20 ns;
input_tb <= "01100101";
wait for 20 ns;
input_tb <= "10000000";
wait for 20 ns;
input_tb <= "00101101";
wait for 20 ns;
input_tb <= "10011010";
wait for 20 ns;
input_tb <= "10100011";
wait for 20 ns;
input_tb <= "10001011";
wait for 20 ns;
input_tb <= "11111001";
wait for 20 ns;
input_tb <= "10101011";
wait for 20 ns;
input_tb <= "01010101";
wait for 20 ns;
input_tb <= "00001101";
wait for 20 ns;
input_tb <= "11101111";
wait for 20 ns;
input_tb <= "10010111";
wait for 20 ns;
input_tb <= "01100110";
wait for 20 ns;
input_tb <= "10010010";
wait for 20 ns;
input_tb <= "01111010";
wait for 20 ns;
input_tb <= "11101011";
wait for 20 ns;
input_tb <= "11001001";
wait for 20 ns;
input_tb <= "10010001";
wait for 20 ns;
input_tb <= "01000001";
wait for 20 ns;
input_tb <= "10000110";
wait for 20 ns;
input_tb <= "01101010";
wait for 20 ns;
input_tb <= "10010110";
wait for 20 ns;
input_tb <= "10110100";
wait for 20 ns;
input_tb <= "11100100";
wait for 20 ns;
input_tb <= "01100101";
wait for 20 ns;
input_tb <= "10100000";
wait for 20 ns;
input_tb <= "11100101";
wait for 20 ns;
input_tb <= "10100011";
wait for 20 ns;
input_tb <= "01110111";
wait for 20 ns;
input_tb <= "11001000";
wait for 20 ns;
input_tb <= "10011010";
wait for 20 ns;
input_tb <= "00111111";
wait for 20 ns;
input_tb <= "10110001";
wait for 20 ns;
input_tb <= "00100100";
wait for 20 ns;
input_tb <= "10100000";
wait for 20 ns;
input_tb <= "00100001";
wait for 20 ns;
input_tb <= "01110100";
wait for 20 ns;
input_tb <= "11101011";
wait for 20 ns;
input_tb <= "01100010";
wait for 20 ns;
input_tb <= "11011000";
wait for 20 ns;
input_tb <= "10011001";
wait for 20 ns;
input_tb <= "11011010";
wait for 20 ns;
input_tb <= "10111010";
wait for 20 ns;
input_tb <= "10100110";
wait for 20 ns;
input_tb <= "11110000";
wait for 20 ns;
input_tb <= "11010110";
wait for 20 ns;
input_tb <= "00000110";
wait for 20 ns;
input_tb <= "00111110";
wait for 20 ns;
input_tb <= "11101100";
wait for 20 ns;
input_tb <= "11010010";
wait for 20 ns;
input_tb <= "01111111";
wait for 20 ns;
input_tb <= "11001100";
wait for 20 ns;
input_tb <= "10011100";
wait for 20 ns;
input_tb <= "11110011";
wait for 20 ns;
input_tb <= "11000110";
wait for 20 ns;
input_tb <= "00110110";
wait for 20 ns;
input_tb <= "11011101";
wait for 20 ns;
input_tb <= "11110010";
wait for 20 ns;
input_tb <= "11000000";
wait for 20 ns;
input_tb <= "10100001";
wait for 20 ns;
input_tb <= "11001111";
wait for 20 ns;
input_tb <= "11000011";
wait for 20 ns;
input_tb <= "10100100";
wait for 20 ns;
input_tb <= "00111000";
wait for 20 ns;
input_tb <= "10000101";
wait for 20 ns;
input_tb <= "01110100";
wait for 20 ns;
input_tb <= "01010010";
wait for 20 ns;
input_tb <= "00101000";
wait for 20 ns;
input_tb <= "00000001";
wait for 20 ns;
input_tb <= "01010111";
wait for 20 ns;
input_tb <= "11100111";
wait for 20 ns;
input_tb <= "11101111";
wait for 20 ns;
input_tb <= "01011111";
wait for 20 ns;
input_tb <= "01100011";
wait for 20 ns;
input_tb <= "10001110";
wait for 20 ns;
input_tb <= "11010111";
wait for 20 ns;
input_tb <= "01010000";
wait for 20 ns;
input_tb <= "11011000";
wait for 20 ns;
input_tb <= "10011001";
wait for 20 ns;
input_tb <= "10111101";
wait for 20 ns;
input_tb <= "11001010";
wait for 20 ns;
input_tb <= "00100010";
wait for 20 ns;
input_tb <= "11010000";
wait for 20 ns;
input_tb <= "00010111";
wait for 20 ns;
input_tb <= "11111110";
wait for 20 ns;
input_tb <= "00000000";
wait for 20 ns;
input_tb <= "00001000";
wait for 20 ns;
input_tb <= "00110110";
wait for 20 ns;
input_tb <= "10001011";
wait for 20 ns;
input_tb <= "11100101";
wait for 20 ns;
input_tb <= "11111000";
wait for 20 ns;
input_tb <= "11001000";
wait for 20 ns;
input_tb <= "11110001";
wait for 20 ns;
input_tb <= "10011111";
wait for 20 ns;
input_tb <= "01001001";
wait for 20 ns;
input_tb <= "10100000";
wait for 20 ns;
input_tb <= "01001000";
wait for 20 ns;
input_tb <= "00110110";
wait for 20 ns;
input_tb <= "11101100";
wait for 20 ns;
input_tb <= "10111010";
wait for 20 ns;
input_tb <= "00110010";
wait for 20 ns;
input_tb <= "00010111";
wait for 20 ns;
input_tb <= "10110000";
wait for 20 ns;
input_tb <= "01111001";
wait for 20 ns;
input_tb <= "00001110";
wait for 20 ns;
input_tb <= "01110001";
wait for 20 ns;
input_tb <= "00010100";
wait for 20 ns;
input_tb <= "00110100";
wait for 20 ns;
input_tb <= "01101110";
wait for 20 ns;
input_tb <= "11100000";
wait for 20 ns;
input_tb <= "01011001";
wait for 20 ns;
input_tb <= "11110001";
wait for 20 ns;
input_tb <= "11001011";
wait for 20 ns;
input_tb <= "01001001";
wait for 20 ns;
input_tb <= "11011100";
wait for 20 ns;
input_tb <= "01110000";
wait for 20 ns;
input_tb <= "01111000";
wait for 20 ns;
input_tb <= "00000101";
wait for 20 ns;
input_tb <= "10100011";
wait for 20 ns;
input_tb <= "01101100";
wait for 20 ns;
input_tb <= "11010101";
wait for 20 ns;
input_tb <= "01000001";
wait for 20 ns;
input_tb <= "00110110";
wait for 20 ns;
input_tb <= "00011101";
wait for 20 ns;
input_tb <= "11000101";
wait for 20 ns;
input_tb <= "10100100";
wait for 20 ns;
input_tb <= "10110000";
wait for 20 ns;
input_tb <= "00000001";
wait for 20 ns;
input_tb <= "01100010";
wait for 20 ns;
input_tb <= "00110011";
wait for 20 ns;
input_tb <= "00010101";
wait for 20 ns;
input_tb <= "11011100";
wait for 20 ns;
input_tb <= "11101111";
wait for 20 ns;
input_tb <= "01110010";
wait for 20 ns;
input_tb <= "11100110";
wait for 20 ns;
input_tb <= "11111110";
wait for 20 ns;
input_tb <= "00001101";
wait for 20 ns;
input_tb <= "11001100";
wait for 20 ns;
input_tb <= "11110011";
wait for 20 ns;
input_tb <= "11000100";
wait for 20 ns;
input_tb <= "00110010";
wait for 20 ns;
input_tb <= "00110101";
wait for 20 ns;
input_tb <= "01110001";
wait for 20 ns;
input_tb <= "01100001";
wait for 20 ns;
input_tb <= "01011000";
wait for 20 ns;
input_tb <= "00001110";
wait for 20 ns;
input_tb <= "01001100";
wait for 20 ns;
input_tb <= "11011110";
wait for 20 ns;
input_tb <= "11110010";
wait for 20 ns;
input_tb <= "01001001";
wait for 20 ns;
input_tb <= "10111111";
wait for 20 ns;
input_tb <= "01100000";
wait for 20 ns;
input_tb <= "00100100";
wait for 20 ns;
input_tb <= "11001101";
wait for 20 ns;
input_tb <= "00100001";
wait for 20 ns;
input_tb <= "10101010";
wait for 20 ns;
input_tb <= "00110011";
wait for 20 ns;
input_tb <= "00011100";
wait for 20 ns;
input_tb <= "00000010";
wait for 20 ns;
input_tb <= "11100010";
wait for 20 ns;
input_tb <= "00111011";
wait for 20 ns;
input_tb <= "00110011";
wait for 20 ns;
input_tb <= "01110110";
wait for 20 ns;
input_tb <= "10011000";
wait for 20 ns;
input_tb <= "00100000";
wait for 20 ns;
input_tb <= "10110010";
wait for 20 ns;
input_tb <= "10110001";
wait for 20 ns;
input_tb <= "00000100";
wait for 20 ns;
input_tb <= "11000110";
wait for 20 ns;
input_tb <= "00111100";
wait for 20 ns;
input_tb <= "11010100";
wait for 20 ns;
input_tb <= "10001111";
wait for 20 ns;
input_tb <= "10000101";
wait for 20 ns;
input_tb <= "00100001";
wait for 20 ns;
input_tb <= "00000111";
wait for 20 ns;
input_tb <= "10010110";
wait for 20 ns;
input_tb <= "11010111";
wait for 20 ns;
input_tb <= "00111010";
wait for 20 ns;
input_tb <= "11001000";
wait for 20 ns;
input_tb <= "01101010";
wait for 20 ns;
input_tb <= "01010100";
wait for 20 ns;
input_tb <= "00010101";
wait for 20 ns;
input_tb <= "10000010";
wait for 20 ns;
input_tb <= "10011011";
wait for 20 ns;
input_tb <= "11100001";
wait for 20 ns;
input_tb <= "01010010";
wait for 20 ns;
input_tb <= "01100010";
wait for 20 ns;
input_tb <= "01110110";
wait for 20 ns;
input_tb <= "00100100";
wait for 20 ns;
input_tb <= "01001101";
wait for 20 ns;
input_tb <= "01100110";
wait for 20 ns;
input_tb <= "11001100";
wait for 20 ns;
input_tb <= "00111011";
wait for 20 ns;
input_tb <= "11111110";
wait for 20 ns;
input_tb <= "10110111";
wait for 20 ns;
input_tb <= "11110101";
wait for 20 ns;
input_tb <= "10101101";
wait for 20 ns;
input_tb <= "00011101";
wait for 20 ns;
input_tb <= "00111000";
wait for 20 ns;
input_tb <= "00010101";
wait;
end process;
end beh;