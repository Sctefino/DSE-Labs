library ieee;
use ieee.std_logic_1164.all;

entity digital_filter is
end digital_filter;

architecture beh of digital_filter is
begin
end beh;